library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
package LED_LUT_pkg is
type array_1d is array (0 to 255) of integer;
constant d2d_LUT : array_1d := (
( 0 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 1 ),
( 2 ),
( 2 ),
( 2 ),
( 2 ),
( 2 ),
( 2 ),
( 2 ),
( 2 ),
( 2 ),
( 3 ),
( 3 ),
( 3 ),
( 3 ),
( 3 ),
( 3 ),
( 3 ),
( 4 ),
( 4 ),
( 4 ),
( 4 ),
( 4 ),
( 4 ),
( 5 ),
( 5 ),
( 5 ),
( 5 ),
( 5 ),
( 6 ),
( 6 ),
( 6 ),
( 6 ),
( 7 ),
( 7 ),
( 7 ),
( 7 ),
( 7 ),
( 8 ),
( 8 ),
( 8 ),
( 9 ),
( 9 ),
( 9 ),
( 9 ),
( 10 ),
( 10 ),
( 10 ),
( 11 ),
( 11 ),
( 11 ),
( 12 ),
( 12 ),
( 12 ),
( 13 ),
( 13 ),
( 13 ),
( 14 ),
( 14 ),
( 14 ),
( 15 ),
( 15 ),
( 16 ),
( 16 ),
( 16 ),
( 17 ),
( 17 ),
( 18 ),
( 18 ),
( 19 ),
( 19 ),
( 19 ),
( 20 ),
( 20 ),
( 21 ),
( 21 ),
( 22 ),
( 22 ),
( 23 ),
( 23 ),
( 24 ),
( 24 ),
( 25 ),
( 26 ),
( 26 ),
( 27 ),
( 27 ),
( 28 ),
( 28 ),
( 29 ),
( 30 ),
( 30 ),
( 31 ),
( 31 ),
( 32 ),
( 33 ),
( 33 ),
( 34 ),
( 35 ),
( 35 ),
( 36 ),
( 37 ),
( 38 ),
( 38 ),
( 39 ),
( 40 ),
( 40 ),
( 41 ),
( 42 ),
( 43 ),
( 44 ),
( 44 ),
( 45 ),
( 46 ),
( 47 ),
( 48 ),
( 48 ),
( 49 ),
( 50 ),
( 51 ),
( 52 ),
( 53 ),
( 54 ),
( 55 ),
( 55 ),
( 56 ),
( 57 ),
( 58 ),
( 59 ),
( 60 ),
( 61 ),
( 62 ),
( 63 ),
( 64 ),
( 65 ),
( 66 ),
( 67 ),
( 68 ),
( 69 ),
( 70 ),
( 71 ),
( 73 ),
( 74 ),
( 75 ),
( 76 ),
( 77 ),
( 78 ),
( 79 ),
( 81 ),
( 82 ),
( 83 ),
( 84 ),
( 85 ),
( 87 ),
( 88 ),
( 89 ),
( 90 ),
( 92 ),
( 93 ),
( 94 ),
( 96 ),
( 97 ),
( 98 ),
( 100 ),
( 101 ),
( 102 ),
( 104 ),
( 105 ),
( 106 ),
( 108 ),
( 109 ),
( 111 ),
( 112 ),
( 114 ),
( 115 ),
( 117 ),
( 118 ),
( 120 ),
( 121 ),
( 123 ),
( 124 ),
( 126 ),
( 128 ),
( 129 ),
( 131 ),
( 132 ),
( 134 ),
( 136 ),
( 137 ),
( 139 ),
( 141 ),
( 143 ),
( 144 ),
( 146 ),
( 148 ),
( 150 ),
( 151 ),
( 153 ),
( 155 ),
( 157 ),
( 159 ),
( 160 ),
( 162 ),
( 164 ),
( 166 ),
( 168 ),
( 170 ),
( 172 ),
( 174 ),
( 176 ),
( 178 ),
( 180 ),
( 182 ),
( 184 ),
( 186 ),
( 188 ),
( 190 ),
( 192 ),
( 194 ),
( 196 ),
( 198 ),
( 201 ),
( 203 ),
( 205 ),
( 207 ),
( 209 ),
( 212 ),
( 214 ),
( 216 ),
( 218 ),
( 221 ),
( 223 ),
( 225 ),
( 228 ),
( 230 ),
( 232 ),
( 235 ),
( 237 ),
( 240 ),
( 242 ),
( 244 ),
( 247 ),
( 249 ),
( 252 ),
( 254 ));
end package LED_LUT_pkg;
