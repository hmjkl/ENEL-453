library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- This is the default LUT_pkg.vhd. It is used for the testbench code (not the
-- RTL). The real LUT_pkg is called "LUT_pkg.vhd"
package LUT_pkg is

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	7381	)	,
(	7366	)	,
(	7352	)	,
(	7338	)	,
(	7323	)	,
(	7309	)	,
(	7294	)	,
(	7280	)	,
(	7266	)	,
(	7252	)	,
(	7237	)	,
(	7223	)	,
(	7209	)	,
(	7195	)	,
(	7181	)	,
(	7167	)	,
(	7152	)	,
(	7138	)	,
(	7124	)	,
(	7110	)	,
(	7096	)	,
(	7082	)	,
(	7068	)	,
(	7055	)	,
(	7041	)	,
(	7027	)	,
(	7013	)	,
(	6999	)	,
(	6985	)	,
(	6972	)	,
(	6958	)	,
(	6944	)	,
(	6930	)	,
(	6917	)	,
(	6903	)	,
(	6889	)	,
(	6876	)	,
(	6862	)	,
(	6849	)	,
(	6835	)	,
(	6822	)	,
(	6808	)	,
(	6795	)	,
(	6781	)	,
(	6768	)	,
(	6754	)	,
(	6741	)	,
(	6728	)	,
(	6714	)	,
(	6701	)	,
(	6688	)	,
(	6675	)	,
(	6661	)	,
(	6648	)	,
(	6635	)	,
(	6622	)	,
(	6609	)	,
(	6596	)	,
(	6583	)	,
(	6569	)	,
(	6556	)	,
(	6543	)	,
(	6530	)	,
(	6517	)	,
(	6505	)	,
(	6492	)	,
(	6479	)	,
(	6466	)	,
(	6453	)	,
(	6440	)	,
(	6427	)	,
(	6415	)	,
(	6402	)	,
(	6389	)	,
(	6376	)	,
(	6364	)	,
(	6351	)	,
(	6338	)	,
(	6326	)	,
(	6313	)	,
(	6300	)	,
(	6288	)	,
(	6275	)	,
(	6263	)	,
(	6250	)	,
(	6238	)	,
(	6225	)	,
(	6213	)	,
(	6201	)	,
(	6188	)	,
(	6176	)	,
(	6163	)	,
(	6151	)	,
(	6139	)	,
(	6127	)	,
(	6114	)	,
(	6102	)	,
(	6090	)	,
(	6078	)	,
(	6066	)	,
(	6053	)	,
(	6041	)	,
(	6029	)	,
(	6017	)	,
(	6005	)	,
(	5993	)	,
(	5981	)	,
(	5969	)	,
(	5957	)	,
(	5945	)	,
(	5933	)	,
(	5921	)	,
(	5910	)	,
(	5898	)	,
(	5886	)	,
(	5874	)	,
(	5862	)	,
(	5850	)	,
(	5839	)	,
(	5827	)	,
(	5815	)	,
(	5804	)	,
(	5792	)	,
(	5780	)	,
(	5769	)	,
(	5757	)	,
(	5746	)	,
(	5734	)	,
(	5722	)	,
(	5711	)	,
(	5699	)	,
(	5688	)	,
(	5677	)	,
(	5665	)	,
(	5654	)	,
(	5642	)	,
(	5631	)	,
(	5620	)	,
(	5608	)	,
(	5597	)	,
(	5586	)	,
(	5574	)	,
(	5563	)	,
(	5552	)	,
(	5541	)	,
(	5530	)	,
(	5518	)	,
(	5507	)	,
(	5496	)	,
(	5485	)	,
(	5474	)	,
(	5463	)	,
(	5452	)	,
(	5441	)	,
(	5430	)	,
(	5419	)	,
(	5408	)	,
(	5397	)	,
(	5386	)	,
(	5375	)	,
(	5364	)	,
(	5354	)	,
(	5343	)	,
(	5332	)	,
(	5321	)	,
(	5310	)	,
(	5300	)	,
(	5289	)	,
(	5278	)	,
(	5268	)	,
(	5257	)	,
(	5246	)	,
(	5236	)	,
(	5225	)	,
(	5215	)	,
(	5204	)	,
(	5193	)	,
(	5183	)	,
(	5172	)	,
(	5162	)	,
(	5151	)	,
(	5141	)	,
(	5131	)	,
(	5120	)	,
(	5110	)	,
(	5099	)	,
(	5089	)	,
(	5079	)	,
(	5068	)	,
(	5058	)	,
(	5048	)	,
(	5038	)	,
(	5027	)	,
(	5017	)	,
(	5007	)	,
(	4997	)	,
(	4987	)	,
(	4977	)	,
(	4967	)	,
(	4956	)	,
(	4946	)	,
(	4936	)	,
(	4926	)	,
(	4916	)	,
(	4906	)	,
(	4896	)	,
(	4886	)	,
(	4876	)	,
(	4867	)	,
(	4857	)	,
(	4847	)	,
(	4837	)	,
(	4827	)	,
(	4817	)	,
(	4807	)	,
(	4798	)	,
(	4788	)	,
(	4778	)	,
(	4768	)	,
(	4759	)	,
(	4749	)	,
(	4739	)	,
(	4730	)	,
(	4720	)	,
(	4711	)	,
(	4701	)	,
(	4691	)	,
(	4682	)	,
(	4672	)	,
(	4663	)	,
(	4653	)	,
(	4644	)	,
(	4634	)	,
(	4625	)	,
(	4615	)	,
(	4606	)	,
(	4597	)	,
(	4587	)	,
(	4578	)	,
(	4569	)	,
(	4559	)	,
(	4550	)	,
(	4541	)	,
(	4532	)	,
(	4522	)	,
(	4513	)	,
(	4504	)	,
(	4495	)	,
(	4486	)	,
(	4476	)	,
(	4467	)	,
(	4458	)	,
(	4449	)	,
(	4440	)	,
(	4431	)	,
(	4422	)	,
(	4413	)	,
(	4404	)	,
(	4395	)	,
(	4386	)	,
(	4377	)	,
(	4368	)	,
(	4359	)	,
(	4350	)	,
(	4341	)	,
(	4333	)	,
(	4324	)	,
(	4315	)	,
(	4306	)	,
(	4297	)	,
(	4288	)	,
(	4280	)	,
(	4271	)	,
(	4262	)	,
(	4254	)	,
(	4245	)	,
(	4236	)	,
(	4228	)	,
(	4219	)	,
(	4210	)	,
(	4202	)	,
(	4193	)	,
(	4185	)	,
(	4176	)	,
(	4168	)	,
(	4159	)	,
(	4151	)	,
(	4142	)	,
(	4134	)	,
(	4125	)	,
(	4117	)	,
(	4108	)	,
(	4100	)	,
(	4092	)	,
(	4083	)	,
(	4075	)	,
(	4067	)	,
(	4058	)	,
(	4050	)	,
(	4042	)	,
(	4034	)	,
(	4025	)	,
(	4017	)	,
(	4009	)	,
(	4001	)	,
(	3993	)	,
(	3984	)	,
(	3976	)	,
(	3968	)	,
(	3960	)	,
(	3952	)	,
(	3944	)	,
(	3936	)	,
(	3928	)	,
(	3920	)	,
(	3912	)	,
(	3904	)	,
(	3896	)	,
(	3888	)	,
(	3880	)	,
(	3872	)	,
(	3864	)	,
(	3856	)	,
(	3848	)	,
(	3841	)	,
(	3833	)	,
(	3825	)	,
(	3817	)	,
(	3809	)	,
(	3802	)	,
(	3794	)	,
(	3786	)	,
(	3778	)	,
(	3771	)	,
(	3763	)	,
(	3755	)	,
(	3748	)	,
(	3740	)	,
(	3732	)	,
(	3725	)	,
(	3717	)	,
(	3710	)	,
(	3702	)	,
(	3694	)	,
(	3687	)	,
(	3679	)	,
(	3672	)	,
(	3664	)	,
(	3657	)	,
(	3650	)	,
(	3642	)	,
(	3635	)	,
(	3627	)	,
(	3620	)	,
(	3613	)	,
(	3605	)	,
(	3598	)	,
(	3591	)	,
(	3583	)	,
(	3576	)	,
(	3569	)	,
(	3561	)	,
(	3554	)	,
(	3547	)	,
(	3540	)	,
(	3533	)	,
(	3525	)	,
(	3518	)	,
(	3511	)	,
(	3504	)	,
(	3497	)	,
(	3490	)	,
(	3483	)	,
(	3476	)	,
(	3468	)	,
(	3461	)	,
(	3454	)	,
(	3447	)	,
(	3440	)	,
(	3433	)	,
(	3426	)	,
(	3419	)	,
(	3413	)	,
(	3406	)	,
(	3399	)	,
(	3392	)	,
(	3385	)	,
(	3378	)	,
(	3371	)	,
(	3364	)	,
(	3358	)	,
(	3351	)	,
(	3344	)	,
(	3337	)	,
(	3330	)	,
(	3324	)	,
(	3317	)	,
(	3310	)	,
(	3304	)	,
(	3297	)	,
(	3290	)	,
(	3284	)	,
(	3277	)	,
(	3270	)	,
(	3264	)	,
(	3257	)	,
(	3251	)	,
(	3244	)	,
(	3237	)	,
(	3231	)	,
(	3224	)	,
(	3218	)	,
(	3211	)	,
(	3205	)	,
(	3198	)	,
(	3192	)	,
(	3185	)	,
(	3179	)	,
(	3173	)	,
(	3166	)	,
(	3160	)	,
(	3154	)	,
(	3147	)	,
(	3141	)	,
(	3135	)	,
(	3128	)	,
(	3122	)	,
(	3116	)	,
(	3109	)	,
(	3103	)	,
(	3097	)	,
(	3091	)	,
(	3084	)	,
(	3078	)	,
(	3072	)	,
(	3066	)	,
(	3060	)	,
(	3054	)	,
(	3047	)	,
(	3041	)	,
(	3035	)	,
(	3029	)	,
(	3023	)	,
(	3017	)	,
(	3011	)	,
(	3005	)	,
(	2999	)	,
(	2993	)	,
(	2987	)	,
(	2981	)	,
(	2975	)	,
(	2969	)	,
(	2963	)	,
(	2957	)	,
(	2951	)	,
(	2945	)	,
(	2939	)	,
(	2934	)	,
(	2928	)	,
(	2922	)	,
(	2916	)	,
(	2910	)	,
(	2904	)	,
(	2899	)	,
(	2893	)	,
(	2887	)	,
(	2881	)	,
(	2876	)	,
(	2870	)	,
(	2864	)	,
(	2859	)	,
(	2853	)	,
(	2847	)	,
(	2842	)	,
(	2836	)	,
(	2830	)	,
(	2825	)	,
(	2819	)	,
(	2813	)	,
(	2808	)	,
(	2802	)	,
(	2797	)	,
(	2791	)	,
(	2786	)	,
(	2780	)	,
(	2775	)	,
(	2769	)	,
(	2764	)	,
(	2758	)	,
(	2753	)	,
(	2747	)	,
(	2742	)	,
(	2736	)	,
(	2731	)	,
(	2726	)	,
(	2720	)	,
(	2715	)	,
(	2710	)	,
(	2704	)	,
(	2699	)	,
(	2694	)	,
(	2688	)	,
(	2683	)	,
(	2678	)	,
(	2673	)	,
(	2667	)	,
(	2662	)	,
(	2657	)	,
(	2652	)	,
(	2646	)	,
(	2641	)	,
(	2636	)	,
(	2631	)	,
(	2626	)	,
(	2621	)	,
(	2615	)	,
(	2610	)	,
(	2605	)	,
(	2600	)	,
(	2595	)	,
(	2590	)	,
(	2585	)	,
(	2580	)	,
(	2575	)	,
(	2570	)	,
(	2565	)	,
(	2560	)	,
(	2555	)	,
(	2550	)	,
(	2545	)	,
(	2540	)	,
(	2535	)	,
(	2530	)	,
(	2525	)	,
(	2520	)	,
(	2515	)	,
(	2511	)	,
(	2506	)	,
(	2501	)	,
(	2496	)	,
(	2491	)	,
(	2486	)	,
(	2482	)	,
(	2477	)	,
(	2472	)	,
(	2467	)	,
(	2463	)	,
(	2458	)	,
(	2453	)	,
(	2448	)	,
(	2444	)	,
(	2439	)	,
(	2434	)	,
(	2430	)	,
(	2425	)	,
(	2420	)	,
(	2416	)	,
(	2411	)	,
(	2406	)	,
(	2402	)	,
(	2397	)	,
(	2393	)	,
(	2388	)	,
(	2383	)	,
(	2379	)	,
(	2374	)	,
(	2370	)	,
(	2365	)	,
(	2361	)	,
(	2356	)	,
(	2352	)	,
(	2347	)	,
(	2343	)	,
(	2338	)	,
(	2334	)	,
(	2330	)	,
(	2325	)	,
(	2321	)	,
(	2316	)	,
(	2312	)	,
(	2308	)	,
(	2303	)	,
(	2299	)	,
(	2295	)	,
(	2290	)	,
(	2286	)	,
(	2282	)	,
(	2277	)	,
(	2273	)	,
(	2269	)	,
(	2264	)	,
(	2260	)	,
(	2256	)	,
(	2252	)	,
(	2247	)	,
(	2243	)	,
(	2239	)	,
(	2235	)	,
(	2231	)	,
(	2227	)	,
(	2222	)	,
(	2218	)	,
(	2214	)	,
(	2210	)	,
(	2206	)	,
(	2202	)	,
(	2198	)	,
(	2194	)	,
(	2189	)	,
(	2185	)	,
(	2181	)	,
(	2177	)	,
(	2173	)	,
(	2169	)	,
(	2165	)	,
(	2161	)	,
(	2157	)	,
(	2153	)	,
(	2149	)	,
(	2145	)	,
(	2141	)	,
(	2137	)	,
(	2134	)	,
(	2130	)	,
(	2126	)	,
(	2122	)	,
(	2118	)	,
(	2114	)	,
(	2110	)	,
(	2106	)	,
(	2102	)	,
(	2099	)	,
(	2095	)	,
(	2091	)	,
(	2087	)	,
(	2083	)	,
(	2080	)	,
(	2076	)	,
(	2072	)	,
(	2068	)	,
(	2064	)	,
(	2061	)	,
(	2057	)	,
(	2053	)	,
(	2050	)	,
(	2046	)	,
(	2042	)	,
(	2039	)	,
(	2035	)	,
(	2031	)	,
(	2028	)	,
(	2024	)	,
(	2020	)	,
(	2017	)	,
(	2013	)	,
(	2009	)	,
(	2006	)	,
(	2002	)	,
(	1999	)	,
(	1995	)	,
(	1991	)	,
(	1988	)	,
(	1984	)	,
(	1981	)	,
(	1977	)	,
(	1974	)	,
(	1970	)	,
(	1967	)	,
(	1963	)	,
(	1960	)	,
(	1956	)	,
(	1953	)	,
(	1950	)	,
(	1946	)	,
(	1943	)	,
(	1939	)	,
(	1936	)	,
(	1932	)	,
(	1929	)	,
(	1926	)	,
(	1922	)	,
(	1919	)	,
(	1916	)	,
(	1912	)	,
(	1909	)	,
(	1906	)	,
(	1902	)	,
(	1899	)	,
(	1896	)	,
(	1892	)	,
(	1889	)	,
(	1886	)	,
(	1882	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1870	)	,
(	1866	)	,
(	1863	)	,
(	1860	)	,
(	1857	)	,
(	1853	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1835	)	,
(	1831	)	,
(	1828	)	,
(	1825	)	,
(	1822	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1804	)	,
(	1801	)	,
(	1798	)	,
(	1795	)	,
(	1792	)	,
(	1789	)	,
(	1786	)	,
(	1783	)	,
(	1780	)	,
(	1777	)	,
(	1774	)	,
(	1771	)	,
(	1768	)	,
(	1765	)	,
(	1762	)	,
(	1759	)	,
(	1756	)	,
(	1753	)	,
(	1750	)	,
(	1747	)	,
(	1744	)	,
(	1742	)	,
(	1739	)	,
(	1736	)	,
(	1733	)	,
(	1730	)	,
(	1727	)	,
(	1724	)	,
(	1722	)	,
(	1719	)	,
(	1716	)	,
(	1713	)	,
(	1710	)	,
(	1708	)	,
(	1705	)	,
(	1702	)	,
(	1699	)	,
(	1697	)	,
(	1694	)	,
(	1691	)	,
(	1688	)	,
(	1686	)	,
(	1683	)	,
(	1680	)	,
(	1678	)	,
(	1675	)	,
(	1672	)	,
(	1670	)	,
(	1667	)	,
(	1664	)	,
(	1662	)	,
(	1659	)	,
(	1656	)	,
(	1654	)	,
(	1651	)	,
(	1648	)	,
(	1646	)	,
(	1643	)	,
(	1641	)	,
(	1638	)	,
(	1636	)	,
(	1633	)	,
(	1630	)	,
(	1628	)	,
(	1625	)	,
(	1623	)	,
(	1620	)	,
(	1618	)	,
(	1615	)	,
(	1613	)	,
(	1610	)	,
(	1608	)	,
(	1605	)	,
(	1603	)	,
(	1600	)	,
(	1598	)	,
(	1595	)	,
(	1593	)	,
(	1590	)	,
(	1588	)	,
(	1586	)	,
(	1583	)	,
(	1581	)	,
(	1578	)	,
(	1576	)	,
(	1574	)	,
(	1571	)	,
(	1569	)	,
(	1566	)	,
(	1564	)	,
(	1562	)	,
(	1559	)	,
(	1557	)	,
(	1555	)	,
(	1552	)	,
(	1550	)	,
(	1548	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1536	)	,
(	1534	)	,
(	1532	)	,
(	1529	)	,
(	1527	)	,
(	1525	)	,
(	1523	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1514	)	,
(	1512	)	,
(	1509	)	,
(	1507	)	,
(	1505	)	,
(	1503	)	,
(	1501	)	,
(	1499	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1431	)	,
(	1429	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1407	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1398	)	,
(	1396	)	,
(	1394	)	,
(	1393	)	,
(	1391	)	,
(	1389	)	,
(	1387	)	,
(	1385	)	,
(	1383	)	,
(	1382	)	,
(	1380	)	,
(	1378	)	,
(	1376	)	,
(	1374	)	,
(	1373	)	,
(	1371	)	,
(	1369	)	,
(	1367	)	,
(	1366	)	,
(	1364	)	,
(	1362	)	,
(	1360	)	,
(	1359	)	,
(	1357	)	,
(	1355	)	,
(	1353	)	,
(	1352	)	,
(	1350	)	,
(	1348	)	,
(	1347	)	,
(	1345	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1338	)	,
(	1337	)	,
(	1335	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1328	)	,
(	1327	)	,
(	1325	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1319	)	,
(	1317	)	,
(	1315	)	,
(	1314	)	,
(	1312	)	,
(	1311	)	,
(	1309	)	,
(	1307	)	,
(	1306	)	,
(	1304	)	,
(	1303	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1295	)	,
(	1294	)	,
(	1292	)	,
(	1290	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1284	)	,
(	1283	)	,
(	1281	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1258	)	,
(	1257	)	,
(	1255	)	,
(	1254	)	,
(	1253	)	,
(	1251	)	,
(	1250	)	,
(	1249	)	,
(	1247	)	,
(	1246	)	,
(	1244	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1235	)	,
(	1234	)	,
(	1232	)	,
(	1231	)	,
(	1230	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1217	)	,
(	1215	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1210	)	,
(	1209	)	,
(	1208	)	,
(	1207	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1202	)	,
(	1200	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1190	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1027	)	,
(	1026	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1015	)	,
(	1014	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1010	)	,
(	1009	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	1000	)	,
(	999	)	,
(	999	)	,
(	998	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	992	)	,
(	991	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	986	)	,
(	985	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	983	)	,
(	982	)	,
(	982	)	,
(	981	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	974	)	,
(	973	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	971	)	,
(	970	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	951	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	362	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	359	)	,
(	358	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	356	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	351	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	349	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	345	)	,
(	345	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	339	)	,
(	339	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	341	)	,
(	341	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	343	)	,
(	343	)	,
(	344	)	,
(	344	)	,
(	345	)	,
(	345	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	347	)	,
(	347	)	,
(	348	)	,
(	348	)	,
(	349	)	,
(	349	)	,
(	350	)	,
(	350	)	,
(	351	)	,
(	351	)	,
(	352	)	,
(	353	)	,
(	353	)	,
(	354	)	,
(	354	)	,
(	355	)	,
(	355	)	,
(	356	)	,
(	356	)	,
(	357	)	,
(	358	)	,
(	358	)	,
(	359	)	,
(	359	)	,
(	360	)	,
(	361	)	,
(	361	)	,
(	362	)	,
(	362	)	,
(	363	)	,
(	364	)	,
(	364	)	,
(	365	)	,
(	366	)	,
(	366	)	,
(	367	)	,
(	368	)	,
(	368	)	,
(	369	)	,
(	370	)	,
(	370	)	,
(	371	)	,
(	372	)	,
(	373	)	,
(	373	)	,
(	374	)	,
(	375	)	,
(	375	)	,
(	376	)	,
(	377	)	,
(	378	)	,
(	378	)	,
(	379	)	,
(	380	)	,
(	381	)	,
(	381	)	,
(	382	)	,
(	383	)	,
(	384	)	,
(	385	)	,
(	385	)	,
(	386	)	,
(	387	)	,
(	388	)	,
(	389	)	,
(	390	)	,
(	390	)	,
(	391	)	,
(	392	)	,
(	393	)	,
(	394	)	,
(	395	)	,
(	396	)	,
(	397	)	,
(	397	)	,
(	398	)	,
(	399	)	,
(	400	)	,
(	401	)	,
(	402	)	,
(	403	)	,
(	404	)	,
(	405	)	,
(	406	)	,
(	407	)	,
(	408	)	,
(	409	)	,
(	410	)	,
(	411	)	,
(	412	)	,
(	413	)	,
(	414	)	,
(	415	)	,
(	416	)	,
(	417	)	,
(	418	)	,
(	419	)	,
(	420	)	,
(	421	)	,
(	422	)	,
(	423	)	,
(	424	)	,
(	425	)	,
(	426	)	,
(	427	)	,
(	428	)	,
(	429	)	,
(	431	)	,
(	432	)	,
(	433	)	,
(	434	)	,
(	435	)	,
(	436	)	,
(	437	)	,
(	438	)	,
(	440	)	,
(	441	)	,
(	442	)	,
(	443	)	,
(	444	)	,
(	446	)	,
(	447	)	,
(	448	)	,
(	449	)	,
(	450	)	,
(	452	)	,
(	453	)	,
(	454	)	,
(	455	)	,
(	457	)	,
(	458	)	,
(	459	)	,
(	460	)	,
(	462	)	,
(	463	)	,
(	464	)	,
(	466	)	,
(	467	)	,
(	468	)	,
(	470	)	,
(	471	)	,
(	472	)	,
(	474	)	,
(	475	)	,
(	476	)	,
(	478	)	,
(	479	)	,
(	480	)	,
(	482	)	,
(	483	)	,
(	485	)	,
(	486	)	,
(	488	)	,
(	489	)	,
(	490	)	,
(	492	)	,
(	493	)	,
(	495	)	,
(	496	)	,
(	498	)	,
(	499	)	,
(	501	)	,
(	502	)	,
(	504	)	,
(	505	)	,
(	507	)	,
(	508	)	,
(	510	)	,
(	511	)	,
(	513	)	,
(	514	)	,
(	516	)	,
(	518	)	,
(	519	)	,
(	521	)	,
(	522	)	,
(	524	)	,
(	526	)	,
(	527	)	,
(	529	)	,
(	531	)	,
(	532	)	,
(	534	)	,
(	535	)	,
(	537	)	,
(	539	)	,
(	540	)	,
(	542	)	,
(	544	)	,
(	546	)	,
(	547	)	,
(	549	)	,
(	551	)	,
(	553	)	,
(	554	)	,
(	556	)	,
(	558	)	,
(	560	)	,
(	561	)	,
(	563	)	,
(	565	)	,
(	567	)	,
(	569	)	,
(	570	)	,
(	572	)	,
(	574	)	,
(	576	)	,
(	578	)	,
(	580	)	,
(	581	)	,
(	583	)	,
(	585	)	,
(	587	)	,
(	589	)	,
(	591	)	,
(	593	)	,
(	595	)	,
(	597	)	,
(	599	)	,
(	601	)	,
(	603	)	,
(	605	)	,
(	607	)	,
(	609	)	,
(	611	)	,
(	613	)	,
(	615	)	,
(	617	)	,
(	619	)	,
(	621	)	,
(	623	)	,
(	625	)	,
(	627	)	,
(	629	)	,
(	631	)	,
(	633	)	,
(	635	)	,
(	637	)	,
(	640	)	,
(	642	)	,
(	644	)	,
(	646	)	,
(	648	)	,
(	650	)	,
(	652	)	,
(	655	)	,
(	657	)	,
(	659	)	,
(	661	)	,
(	663	)	,
(	666	)	,
(	668	)	,
(	670	)	,
(	672	)	,
(	675	)	,
(	677	)	,
(	679	)	,
(	682	)	,
(	684	)	,
(	686	)	,
(	688	)	,
(	691	)	,
(	693	)	,
(	696	)	,
(	698	)	,
(	700	)	,
(	703	)	,
(	705	)	,
(	707	)	,
(	710	)	,
(	712	)	,
(	715	)	,
(	717	)	,
(	720	)	,
(	722	)	,
(	724	)	,
(	727	)	,
(	729	)	,
(	732	)	,
(	734	)	,
(	737	)	,
(	739	)	,
(	742	)	,
(	744	)	,
(	747	)	,
(	750	)	,
(	752	)	,
(	755	)	,
(	757	)	,
(	760	)	,
(	763	)	,
(	765	)	,
(	768	)	,
(	770	)	,
(	773	)	,
(	776	)	,
(	778	)	,
(	781	)	,
(	784	)	,
(	786	)	,
(	789	)	,
(	792	)	,
(	795	)	,
(	797	)	,
(	800	)	,
(	803	)	,
(	806	)	,
(	808	)	,
(	811	)	,
(	814	)	,
(	817	)	,
(	820	)	,
(	822	)	,
(	825	)	,
(	828	)	,
(	831	)	,
(	834	)	,
(	837	)	,
(	840	)	,
(	842	)	,
(	845	)	,
(	848	)	,
(	851	)	,
(	854	)	,
(	857	)	,
(	860	)	,
(	863	)	,
(	866	)	,
(	869	)	,
(	872	)	,
(	875	)	,
(	878	)	,
(	881	)	,
(	884	)	,
(	887	)	,
(	890	)	,
(	893	)	,
(	896	)	,
(	899	)	,
(	903	)	,
(	906	)	,
(	909	)	,
(	912	)	,
(	915	)	,
(	918	)	,
(	921	)	,
(	925	)	,
(	928	)	,
(	931	)	,
(	934	)	,
(	937	)	,
(	941	)	,
(	944	)	,
(	947	)	,
(	950	)	,
(	954	)	,
(	957	)	,
(	960	)	,
(	964	)	,
(	967	)	,
(	970	)	,
(	974	)	,
(	977	)	,
(	980	)	,
(	984	)	,
(	987	)	,
(	991	)	,
(	994	)	,
(	997	)	,
(	1001	)	,
(	1004	)	,
(	1008	)	,
(	1011	)	,
(	1015	)	,
(	1018	)	,
(	1022	)	,
(	1025	)	,
(	1029	)	,
(	1032	)	,
(	1036	)	,
(	1039	)	,
(	1043	)	,
(	1047	)	,
(	1050	)	,
(	1054	)	,
(	1057	)	,
(	1061	)	,
(	1065	)	,
(	1068	)	,
(	1072	)	,
(	1076	)	,
(	1079	)	,
(	1083	)	,
(	1087	)	,
(	1091	)	,
(	1094	)	,
(	1098	)	,
(	1102	)	,
(	1106	)	,
(	1109	)	,
(	1113	)	,
(	1117	)	,
(	1121	)	,
(	1125	)	,
(	1128	)	,
(	1132	)	,
(	1136	)	,
(	1140	)	,
(	1144	)	,
(	1148	)	,
(	1152	)	,
(	1156	)	,
(	1160	)	,
(	1164	)	,
(	1168	)	,
(	1172	)	,
(	1176	)	,
(	1180	)	,
(	1184	)	,
(	1188	)	,
(	1192	)	,
(	1196	)	,
(	1200	)	,
(	1204	)	,
(	1208	)	,
(	1212	)	,
(	1216	)	,
(	1220	)	,
(	1224	)	,
(	1228	)	,
(	1233	)	,
(	1237	)	,
(	1241	)	,
(	1245	)	,
(	1249	)	,
(	1254	)	,
(	1258	)	,
(	1262	)	,
(	1266	)	,
(	1271	)	,
(	1275	)	,
(	1279	)	,
(	1284	)	,
(	1288	)	,
(	1292	)	,
(	1297	)	,
(	1301	)	,
(	1305	)	,
(	1310	)	,
(	1314	)	,
(	1319	)	,
(	1323	)	,
(	1327	)	,
(	1332	)	,
(	1336	)	,
(	1341	)	,
(	1345	)	,
(	1350	)	,
(	1354	)	,
(	1359	)	,
(	1363	)	,
(	1368	)	,
(	1373	)	,
(	1377	)	,
(	1382	)	,
(	1386	)	,
(	1391	)	,
(	1396	)	,
(	1400	)	,
(	1405	)	,
(	1410	)	,
(	1414	)	,
(	1419	)	,
(	1424	)	,
(	1428	)	,
(	1433	)	,
(	1438	)	,
(	1443	)	,
(	1448	)	,
(	1452	)	,
(	1457	)	,
(	1462	)	,
(	1467	)	,
(	1472	)	,
(	1477	)	,
(	1481	)	,
(	1486	)	,
(	1491	)	,
(	1496	)	,
(	1501	)	,
(	1506	)	,
(	1511	)	,
(	1516	)	,
(	1521	)	,
(	1526	)	,
(	1531	)	,
(	1536	)	,
(	1541	)	,
(	1546	)	,
(	1551	)	,
(	1556	)	,
(	1561	)	,
(	1567	)	,
(	1572	)	,
(	1577	)	,
(	1582	)	,
(	1587	)	,
(	1592	)	,
(	1597	)	,
(	1603	)	,
(	1608	)	,
(	1613	)	,
(	1618	)	,
(	1624	)	,
(	1629	)	,
(	1634	)	,
(	1640	)	,
(	1645	)	,
(	1650	)	,
(	1656	)	,
(	1661	)	,
(	1666	)	,
(	1672	)	,
(	1677	)	,
(	1683	)	,
(	1688	)	,
(	1694	)	,
(	1699	)	,
(	1705	)	,
(	1710	)	,
(	1716	)	,
(	1721	)	,
(	1727	)	,
(	1732	)	,
(	1738	)	,
(	1743	)	,
(	1749	)	,
(	1755	)	,
(	1760	)	,
(	1766	)	,
(	1772	)	,
(	1777	)	,
(	1783	)	,
(	1789	)	,
(	1794	)	,
(	1800	)	,
(	1806	)	,
(	1812	)	,
(	1817	)	,
(	1823	)	,
(	1829	)	,
(	1835	)	,
(	1841	)	,
(	1847	)	,
(	1852	)	,
(	1858	)	,
(	1864	)	,
(	1870	)	,
(	1876	)	,
(	1882	)	,
(	1888	)	,
(	1894	)	,
(	1900	)	,
(	1906	)	,
(	1912	)	,
(	1918	)	,
(	1924	)	,
(	1930	)	,
(	1936	)	,
(	1942	)	,
(	1948	)	,
(	1955	)	,
(	1961	)	,
(	1967	)	,
(	1973	)	,
(	1979	)	,
(	1986	)	,
(	1992	)	,
(	1998	)	,
(	2004	)	,
(	2011	)	,
(	2017	)	,
(	2023	)	,
(	2029	)	,
(	2036	)	,
(	2042	)	,
(	2049	)	,
(	2055	)	,
(	2061	)	,
(	2068	)	,
(	2074	)	,
(	2081	)	,
(	2087	)	,
(	2094	)	,
(	2100	)	,
(	2107	)	,
(	2113	)	,
(	2120	)	,
(	2126	)	,
(	2133	)	,
(	2139	)	,
(	2146	)	,
(	2153	)	,
(	2159	)	,
(	2166	)	,
(	2173	)	,
(	2179	)	,
(	2186	)	,
(	2193	)	,
(	2200	)	,
(	2206	)	,
(	2213	)	,
(	2220	)	,
(	2227	)	,
(	2233	)	,
(	2240	)	,
(	2247	)	,
(	2254	)	,
(	2261	)	,
(	2268	)	,
(	2275	)	,
(	2282	)	,
(	2289	)	,
(	2296	)	,
(	2303	)	,
(	2310	)	,
(	2317	)	,
(	2324	)	,
(	2331	)	,
(	2338	)	,
(	2345	)	,
(	2352	)	,
(	2359	)	,
(	2366	)	,
(	2374	)	,
(	2381	)	,
(	2388	)	,
(	2395	)	,
(	2402	)	,
(	2410	)	,
(	2417	)	,
(	2424	)	,
(	2431	)	,
(	2439	)	,
(	2446	)	,
(	2453	)	,
(	2461	)	,
(	2468	)	,
(	2476	)	,
(	2483	)	,
(	2490	)	,
(	2498	)	,
(	2505	)	,
(	2513	)	,
(	2520	)	,
(	2528	)	,
(	2535	)	,
(	2543	)	,
(	2551	)	,
(	2558	)	,
(	2566	)	,
(	2573	)	,
(	2581	)	,
(	2589	)	,
(	2596	)	,
(	2604	)	,
(	2612	)	,
(	2620	)	,
(	2627	)	,
(	2635	)	,
(	2643	)	,
(	2651	)	,
(	2658	)	,
(	2666	)	,
(	2674	)	,
(	2682	)	,
(	2690	)	,
(	2698	)	,
(	2706	)	,
(	2714	)	,
(	2722	)	,
(	2730	)	,
(	2738	)	,
(	2746	)	,
(	2754	)	,
(	2762	)	,
(	2770	)	,
(	2778	)	,
(	2786	)	,
(	2794	)	,
(	2802	)	,
(	2811	)	,
(	2819	)	,
(	2827	)	,
(	2835	)	,
(	2843	)	,
(	2852	)	,
(	2860	)	,
(	2868	)	,
(	2877	)	,
(	2885	)	,
(	2893	)	,
(	2902	)	,
(	2910	)	,
(	2919	)	,
(	2927	)	,
(	2935	)	,
(	2944	)	,
(	2952	)	,
(	2961	)	,
(	2969	)	,
(	2978	)	,
(	2987	)	,
(	2995	)	,
(	3004	)	,
(	3012	)	,
(	3021	)	,
(	3030	)	,
(	3038	)	,
(	3047	)	,
(	3056	)	,
(	3064	)	,
(	3073	)	,
(	3082	)	,
(	3091	)	,
(	3100	)	,
(	3108	)	,
(	3117	)	,
(	3126	)	,
(	3135	)	,
(	3144	)	,
(	3153	)	,
(	3162	)	,
(	3171	)	,
(	3180	)	,
(	3189	)	,
(	3198	)	,
(	3207	)	,
(	3216	)	,
(	3225	)	,
(	3234	)	,
(	3243	)	,
(	3252	)	,
(	3261	)	,
(	3271	)	,
(	3280	)	,
(	3289	)	,
(	3298	)	,
(	3308	)	,
(	3317	)	,
(	3326	)	,
(	3335	)	,
(	3345	)	,
(	3354	)	,
(	3364	)	,
(	3373	)	,
(	3382	)	,
(	3392	)	,
(	3401	)	,
(	3411	)	,
(	3420	)	,
(	3430	)	,
(	3439	)	,
(	3449	)	,
(	3458	)	,
(	3468	)	,
(	3478	)	,
(	3487	)	,
(	3497	)	,
(	3507	)	,
(	3516	)	,
(	3526	)	,
(	3536	)	,
(	3546	)	,
(	3555	)	,
(	3565	)	,
(	3575	)	,
(	3585	)	,
(	3595	)	,
(	3605	)	,
(	3615	)	,
(	3624	)	,
(	3634	)	,
(	3644	)	,
(	3654	)	,
(	3664	)	,
(	3674	)	,
(	3684	)	,
(	3695	)	,
(	3705	)	,
(	3715	)	,
(	3725	)	,
(	3735	)	,
(	3745	)	,
(	3755	)	,
(	3766	)	,
(	3776	)	,
(	3786	)	,
(	3796	)	,
(	3807	)	,
(	3817	)	,
(	3827	)	,
(	3838	)	,
(	3848	)	,
(	3859	)	,
(	3869	)	,
(	3879	)	,
(	3890	)	,
(	3900	)	,
(	3911	)	,
(	3922	)	,
(	3932	)	,
(	3943	)	,
(	3953	)	,
(	3964	)	,
(	3975	)	,
(	3985	)	,
(	3996	)	,
(	4007	)	,
(	4017	)	,
(	4028	)	,
(	4039	)	,
(	4050	)	,
(	4060	)	,
(	4071	)	,
(	4082	)	,
(	4093	)	,
(	4104	)	,
(	4115	)	,
(	4126	)	,
(	4137	)	,
(	4148	)	,
(	4159	)	,
(	4170	)	,
(	4181	)	,
(	4192	)	,
(	4203	)	,
(	4214	)	,
(	4225	)	,
(	4237	)	,
(	4248	)	,
(	4259	)	,
(	4270	)	,
(	4282	)	,
(	4293	)	,
(	4304	)	,
(	4315	)	,
(	4327	)	,
(	4338	)	,
(	4350	)	,
(	4361	)	,
(	4372	)	,
(	4384	)	,
(	4395	)	,
(	4407	)	,
(	4418	)	,
(	4430	)	,
(	4442	)	,
(	4453	)	,
(	4465	)	,
(	4476	)	,
(	4488	)	,
(	4500	)	,
(	4512	)	,
(	4523	)	,
(	4535	)	,
(	4547	)	,
(	4559	)	,
(	4570	)	,
(	4582	)	,
(	4594	)	,
(	4606	)	,
(	4618	)	,
(	4630	)	,
(	4642	)	,
(	4654	)	,
(	4666	)	,
(	4678	)	,
(	4690	)	,
(	4702	)	,
(	4714	)	,
(	4726	)	,
(	4738	)	,
(	4751	)	,
(	4763	)	,
(	4775	)	,
(	4787	)	,
(	4800	)	,
(	4812	)	,
(	4824	)	,
(	4837	)	,
(	4849	)	,
(	4861	)	,
(	4874	)	,
(	4886	)	,
(	4899	)	,
(	4911	)	,
(	4924	)	,
(	4936	)	,
(	4949	)	,
(	4961	)	,
(	4974	)	,
(	4987	)	,
(	4999	)	,
(	5012	)	,
(	5025	)	,
(	5037	)	,
(	5050	)	,
(	5063	)	,
(	5076	)	,
(	5088	)	,
(	5101	)	,
(	5114	)	,
(	5127	)	,
(	5140	)	,
(	5153	)	,
(	5166	)	,
(	5179	)	,
(	5192	)	,
(	5205	)	,
(	5218	)	,
(	5231	)	,
(	5244	)	,
(	5257	)	,
(	5270	)	,
(	5284	)	,
(	5297	)	,
(	5310	)	,
(	5323	)	,
(	5337	)	,
(	5350	)	,
(	5363	)	,
(	5377	)	,
(	5390	)	,
(	5403	)	,
(	5417	)	,
(	5430	)	,
(	5444	)	,
(	5457	)	,
(	5471	)	,
(	5484	)	,
(	5498	)	,
(	5512	)	,
(	5525	)	,
(	5539	)	,
(	5553	)	,
(	5566	)	,
(	5580	)	,
(	5594	)	,
(	5608	)	,
(	5621	)	,
(	5635	)	,
(	5649	)	,
(	5663	)	,
(	5677	)	,
(	5691	)	,
(	5705	)	,
(	5719	)	,
(	5733	)	,
(	5747	)	,
(	5761	)	,
(	5775	)	,
(	5789	)	,
(	5803	)	,
(	5817	)	,
(	5832	)	,
(	5846	)	,
(	5860	)	,
(	5874	)	,
(	5889	)	,
(	5903	)	,
(	5917	)	,
(	5932	)	,
(	5946	)	,
(	5961	)	,
(	5975	)	,
(	5989	)	,
(	6004	)	,
(	6018	)	,
(	6033	)	,
(	6048	)	,
(	6062	)	,
(	6077	)	,
(	6092	)	,
(	6106	)	,
(	6121	)	,
(	6136	)	,
(	6150	)	,
(	6165	)	,
(	6180	)	,
(	6195	)	,
(	6210	)	,
(	6225	)	,
(	6240	)	,
(	6255	)	,
(	6270	)	,
(	6285	)	,
(	6300	)	,
(	6315	)	,
(	6330	)	,
(	6345	)	,
(	6360	)	,
(	6375	)	,
(	6390	)	,
(	6406	)	,
(	6421	)	,
(	6436	)	,
(	6451	)	,
(	6467	)	,
(	6482	)	,
(	6497	)	,
(	6513	)	,
(	6528	)	,
(	6544	)	,
(	6559	)	,
(	6575	)	,
(	6590	)	,
(	6606	)	,
(	6622	)	,
(	6637	)	,
(	6653	)	,
(	6668	)	,
(	6684	)	,
(	6700	)	,
(	6716	)	,
(	6732	)	,
(	6747	)	,
(	6763	)	,
(	6779	)	,
(	6795	)	,
(	6811	)	,
(	6827	)	,
(	6843	)	,
(	6859	)	,
(	6875	)	,
(	6891	)	,
(	6907	)	,
(	6923	)	,
(	6939	)	,
(	6956	)	,
(	6972	)	,
(	6988	)	,
(	7004	)	,
(	7021	)	,
(	7037	)	,
(	7053	)	,
(	7070	)	,
(	7086	)	,
(	7102	)	,
(	7119	)	,
(	7135	)	,
(	7152	)	,
(	7168	)	,
(	7185	)	,
(	7202	)	,
(	7218	)	,
(	7235	)	,
(	7252	)	,
(	7268	)	,
(	7285	)	,
(	7302	)	,
(	7319	)	,
(	7335	)	,
(	7352	)	,
(	7369	)	,
(	7386	)	,
(	7403	)	,
(	7420	)	,
(	7437	)	,
(	7454	)	,
(	7471	)	,
(	7488	)	,
(	7505	)	,
(	7523	)	,
(	7540	)	,
(	7557	)	,
(	7574	)	,
(	7591	)	,
(	7609	)	,
(	7626	)	,
(	7643	)	,
(	7661	)	,
(	7678	)	,
(	7696	)	,
(	7713	)	,
(	7731	)	,
(	7748	)	,
(	7766	)	,
(	7783	)	,
(	7801	)	,
(	7819	)	,
(	7836	)	,
(	7854	)	,
(	7872	)	,
(	7889	)	,
(	7907	)	,
(	7925	)	,
(	7943	)	,
(	7961	)	,
(	7979	)	,
(	7997	)	,
(	8015	)	,
(	8033	)	,
(	8051	)	,
(	8069	)	,
(	8087	)	,
(	8105	)	,
(	8123	)	,
(	8141	)	,
(	8159	)	,
(	8178	)	,
(	8196	)	,
(	8214	)	,
(	8233	)	,
(	8251	)	,
(	8269	)	,
(	8288	)	,
(	8306	)	,
(	8325	)	,
(	8343	)	,
(	8362	)	,
(	8380	)	,
(	8399	)	,
(	8418	)	,
(	8436	)	,
(	8455	)	,
(	8474	)	,
(	8493	)	,
(	8511	)	,
(	8530	)	,
(	8549	)	,
(	8568	)	,
(	8587	)	,
(	8606	)	,
(	8625	)	,
(	8644	)	,
(	8663	)	,
(	8682	)	,
(	8701	)	,
(	8720	)	,
(	8739	)	,
(	8758	)	,
(	8778	)	,
(	8797	)	,
(	8816	)	,
(	8835	)	,
(	8855	)	,
(	8874	)	,
(	8894	)	,
(	8913	)	,
(	8933	)	,
(	8952	)	,
(	8972	)	,
(	8991	)	,
(	9011	)	,
(	9030	)	,
(	9050	)	,
(	9070	)	,
(	9089	)	,
(	9109	)	,
(	9129	)	,
(	9149	)	,
(	9169	)	,
(	9189	)	,
(	9209	)	,
(	9228	)	,
(	9248	)	,
(	9268	)	,
(	9289	)	,
(	9309	)	,
(	9329	)	,
(	9349	)	,
(	9369	)	,
(	9389	)	,
(	9409	)	,
(	9430	)	,
(	9450	)	,
(	9470	)	,
(	9491	)	,
(	9511	)	,
(	9532	)	,
(	9552	)	,
(	9573	)	,
(	9593	)	,
(	9614	)	,
(	9634	)	,
(	9655	)	,
(	9676	)	,
(	9696	)	,
(	9717	)	,
(	9738	)	,
(	9758	)	,
(	9779	)	,
(	9800	)	,
(	9821	)	,
(	9842	)	,
(	9863	)	,
(	9884	)	,
(	9905	)	,
(	9926	)	,
(	9947	)	,
(	9968	)	,
(	9989	)	,
(	10011	)	,
(	10032	)	,
(	10053	)	,
(	10074	)	,
(	10096	)	,
(	10117	)	,
(	10138	)	,
(	10160	)	,
(	10181	)	,
(	10203	)	,
(	10224	)	,
(	10246	)	,
(	10267	)	,
(	10289	)	,
(	10311	)	,
(	10332	)	,
(	10354	)	,
(	10376	)	,
(	10398	)	,
(	10419	)	,
(	10441	)	,
(	10463	)	,
(	10485	)	,
(	10507	)	,
(	10529	)	,
(	10551	)	,
(	10573	)	,
(	10595	)	,
(	10617	)	,
(	10639	)	,
(	10662	)	,
(	10684	)	,
(	10706	)	,
(	10728	)	,
(	10751	)	,
(	10773	)	,
(	10796	)	,
(	10818	)	,
(	10840	)	,
(	10863	)	,
(	10885	)	,
(	10908	)	,
(	10931	)	,
(	10953	)	,
(	10976	)	,
(	10999	)	,
(	11021	)	,
(	11044	)	,
(	11067	)	,
(	11090	)	,
(	11113	)	,
(	11136	)	,
(	11159	)	,
(	11182	)	,
(	11205	)	,
(	11228	)	,
(	11251	)	,
(	11274	)	,
(	11297	)	,
(	11320	)	,
(	11343	)	,
(	11367	)	,
(	11390	)	,
(	11413	)	,
(	11437	)	,
(	11460	)	,
(	11484	)	,
(	11507	)	,
(	11531	)	,
(	11554	)	,
(	11578	)	,
(	11601	)	,
(	11625	)	,
(	11649	)	,
(	11672	)	,
(	11696	)	,
(	11720	)	,
(	11744	)	,
(	11768	)	,
(	11792	)	,
(	11816	)	,
(	11840	)	,
(	11864	)	,
(	11888	)	,
(	11912	)	,
(	11936	)	,
(	11960	)	,
(	11984	)	,
(	12008	)	,
(	12033	)	,
(	12057	)	,
(	12081	)	,
(	12106	)	,
(	12130	)	,
(	12155	)	,
(	12179	)	,
(	12204	)	,
(	12228	)	,
(	12253	)	,
(	12277	)	,
(	12302	)	,
(	12327	)	,
(	12351	)	,
(	12376	)	,
(	12401	)	,
(	12426	)	,
(	12451	)	,
(	12476	)	,
(	12501	)	,
(	12526	)	,
(	12551	)	,
(	12576	)	,
(	12601	)	,
(	12626	)	,
(	12651	)	,
(	12676	)	,
(	12702	)	,
(	12727	)	,
(	12752	)	,
(	12778	)	,
(	12803	)	,
(	12828	)	,
(	12854	)	,
(	12879	)	,
(	12905	)	,
(	12931	)	,
(	12956	)	,
(	12982	)	,
(	13008	)	,
(	13033	)	,
(	13059	)	,
(	13085	)	,
(	13111	)	,
(	13137	)	,
(	13163	)	,
(	13189	)	,
(	13215	)	,
(	13241	)	,
(	13267	)	,
(	13293	)	,
(	13319	)	,
(	13345	)	,
(	13371	)	,
(	13398	)	,
(	13424	)	,
(	13450	)	,
(	13477	)	,
(	13503	)	,
(	13529	)	,
(	13556	)	,
(	13583	)	,
(	13609	)	,
(	13636	)	,
(	13662	)	,
(	13689	)	,
(	13716	)	,
(	13743	)	,
(	13769	)	,
(	13796	)	,
(	13823	)	,
(	13850	)	,
(	13877	)	,
(	13904	)	,
(	13931	)	,
(	13958	)	,
(	13985	)	,
(	14012	)	,
(	14039	)	,
(	14067	)	,
(	14094	)	,
(	14121	)	,
(	14149	)	,
(	14176	)	,
(	14203	)	,
(	14231	)	,
(	14258	)	,
(	14286	)	,
(	14314	)	,
(	14341	)	,
(	14369	)	,
(	14396	)	,
(	14424	)	,
(	14452	)	,
(	14480	)	,
(	14508	)	,
(	14536	)	,
(	14563	)	,
(	14591	)	,
(	14619	)	,
(	14648	)	,
(	14676	)	,
(	14704	)	,
(	14732	)	,
(	14760	)	,
(	14788	)	,
(	14817	)	,
(	14845	)	,
(	14873	)	,
(	14902	)	,
(	14930	)	,
(	14959	)	,
(	14987	)	,
(	15016	)	,
(	15044	)	,
(	15073	)	,
(	15102	)	,
(	15130	)	,
(	15159	)	,
(	15188	)	,
(	15217	)	,
(	15246	)	,
(	15275	)	,
(	15304	)	,
(	15333	)	,
(	15362	)	,
(	15391	)	,
(	15420	)	,
(	15449	)	,
(	15478	)	,
(	15508	)	,
(	15537	)	,
(	15566	)	,
(	15596	)	,
(	15625	)	,
(	15655	)	,
(	15684	)	,
(	15714	)	,
(	15743	)	,
(	15773	)	,
(	15802	)	,
(	15832	)	,
(	15862	)	,
(	15892	)	,
(	15922	)	,
(	15951	)	,
(	15981	)	,
(	16011	)	,
(	16041	)	,
(	16071	)	,
(	16101	)	,
(	16132	)
);


end package LUT_pkg;
