library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
package LED_LUT_pkg is
type array_1d is array (0 to 255) of integer;
constant d2d_LUT : array_1d := (
( 23 ),
( 22 ),
( 22 ),
( 21 ),
( 21 ),
( 20 ),
( 20 ),
( 20 ),
( 19 ),
( 19 ),
( 18 ),
( 18 ),
( 18 ),
( 17 ),
( 17 ),
( 17 ),
( 17 ),
( 16 ),
( 16 ),
( 16 ),
( 16 ),
( 16 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 14 ),
( 14 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 15 ),
( 16 ),
( 16 ),
( 16 ),
( 16 ),
( 16 ),
( 17 ),
( 17 ),
( 17 ),
( 18 ),
( 18 ),
( 18 ),
( 18 ),
( 19 ),
( 19 ),
( 19 ),
( 20 ),
( 20 ),
( 21 ),
( 21 ),
( 21 ),
( 22 ),
( 22 ),
( 23 ),
( 23 ),
( 24 ),
( 24 ),
( 25 ),
( 25 ),
( 26 ),
( 26 ),
( 27 ),
( 27 ),
( 28 ),
( 29 ),
( 29 ),
( 30 ),
( 30 ),
( 31 ),
( 32 ),
( 32 ),
( 33 ),
( 34 ),
( 34 ),
( 35 ),
( 36 ),
( 37 ),
( 37 ),
( 38 ),
( 39 ),
( 40 ),
( 40 ),
( 41 ),
( 42 ),
( 43 ),
( 43 ),
( 44 ),
( 45 ),
( 46 ),
( 47 ),
( 48 ),
( 48 ),
( 49 ),
( 50 ),
( 51 ),
( 52 ),
( 53 ),
( 54 ),
( 55 ),
( 56 ),
( 57 ),
( 57 ),
( 58 ),
( 59 ),
( 60 ),
( 61 ),
( 62 ),
( 63 ),
( 64 ),
( 65 ),
( 66 ),
( 67 ),
( 68 ),
( 69 ),
( 70 ),
( 71 ),
( 72 ),
( 74 ),
( 75 ),
( 76 ),
( 77 ),
( 78 ),
( 79 ),
( 80 ),
( 81 ),
( 82 ),
( 83 ),
( 84 ),
( 86 ),
( 87 ),
( 88 ),
( 89 ),
( 90 ),
( 91 ),
( 92 ),
( 94 ),
( 95 ),
( 96 ),
( 97 ),
( 98 ),
( 99 ),
( 101 ),
( 102 ),
( 103 ),
( 104 ),
( 105 ),
( 107 ),
( 108 ),
( 109 ),
( 110 ),
( 112 ),
( 113 ),
( 114 ),
( 115 ),
( 116 ),
( 118 ),
( 119 ),
( 120 ),
( 121 ),
( 123 ),
( 124 ),
( 125 ),
( 126 ),
( 128 ),
( 129 ),
( 130 ),
( 132 ),
( 133 ),
( 134 ),
( 135 ),
( 137 ),
( 138 ),
( 139 ),
( 141 ),
( 142 ),
( 143 ),
( 144 ),
( 146 ),
( 147 ),
( 148 ),
( 150 ),
( 151 ),
( 152 ),
( 154 ),
( 155 ),
( 156 ),
( 157 ),
( 159 ),
( 160 ),
( 161 ),
( 163 ),
( 164 ),
( 165 ),
( 167 ),
( 168 ),
( 169 ),
( 171 ),
( 172 ),
( 173 ),
( 174 ),
( 176 ),
( 177 ),
( 178 ),
( 180 ),
( 181 ),
( 182 ),
( 184 ),
( 185 ),
( 186 ),
( 187 ),
( 189 ),
( 190 ),
( 191 ),
( 193 ),
( 194 ),
( 195 ),
( 197 ),
( 198 ),
( 199 ),
( 200 ),
( 202 ),
( 203 ),
( 204 ),
( 205 ),
( 207 ),
( 208 ),
( 209 ),
( 211 ),
( 212 ),
( 213 ),
( 214 ),
( 216 ),
( 217 ),
( 218 ),
( 219 ),
( 220 ),
( 222 ),
( 223 ),
( 224 ),
( 225 ),
( 227 ),
( 228 ));
end package LED_LUT_pkg;
